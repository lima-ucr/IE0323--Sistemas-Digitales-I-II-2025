module add_sub (
    input [3:0] A,
    input [3:0] B,
    input sum_notsub,
    output reg overflow,
    output reg [3:0] result
);
    
endmodule