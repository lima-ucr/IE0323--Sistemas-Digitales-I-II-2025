module bin_2_seg (
    input [3:0] binary,
    output reg [7:0] segments
);
    
endmodule