module res_to_sign_mag (
    input [3:0] result,
    output reg sign,
    output reg [3:0] magnitude
);
    
endmodule