module mux2x1_param #(
    parameter WIDTH = 8
) (
    input [WIDTH-1:0] D0,
    input [WIDTH-1:0] D1,
    input sel,
    output reg [WIDTH-1:0] Y
);
    
endmodule