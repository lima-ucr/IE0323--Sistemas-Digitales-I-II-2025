module sign_2_seg (
    input sign,
    output reg [7:0] seg
);
    
endmodule